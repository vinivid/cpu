library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity control_unit is
    port (
        instruction : in STD_LOGIC_VECTOR (7 downto 0)
    );
end entity control_unit;

architecture Behaviour of control_unit is
    
begin
    
    
    
end architecture Behaviour;