library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity decoder is
    port (
        
    );
end entity decoder;

architecture Behaviour of decoder is
    
begin
    
    
    
end architecture Behaviour;